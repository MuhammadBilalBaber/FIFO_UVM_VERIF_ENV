package fifo_package;
  `include "uvm_macros.svh"
   import uvm_pkg::*;
   `include "fifo_seq_item.sv"
   `include "fifo_sequence.sv"
   `include "fifo_read_sequence.sv"
   `include "fifo_sequencer.sv"
   `include "fifo_read_sequencer.sv"
   `include "fifo_virtual_sequencer.sv"
   `include "fifo_virtual_sequence.sv"
   `include "fifo_driver.sv"
   `include "fifo_read_driver.sv"
   `include "fifo_monitor.sv"
   `include "fifo_read_monitor.sv"
   `include "fifo_agent.sv"
   `include "fifo_read_agent.sv"
   `include "fifo_environment.sv"
   `include "fifo_test.sv"

endpackage : fifo_package